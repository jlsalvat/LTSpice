* HCMOS Subcircuit and Primitive Elements Library
* HC_TSLOW.CIR
* Slow Process Corner
* Standard Logic Product Group
* Philips Semiconductors
*
* Version Date       By   Remarks
* ---------------------------------------------------------------------
*    1.05 10/27/2005 RRV  Updated HC/T04 and HCU04 models
*    1.04 09/22/2003 RM   Active High Enable for SWI2 and SWI2T
*
************************************************
*          SLOW N-Channel Transistor           *
*            UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family         *
*                10-Jan.-1995                  *
************************************************
.Model MHCNES NMOS
+LEVEL = 3
+KP    = 41.0E-6
+VTO   = 0.92
+TOX   = 54.0E-9
+NSUB  = 2.0E15
+GAMMA = 1.14
+PHI   = 0.65
+VMAX  = 175E3
+RS    = 50
+RD    = 50
+XJ    = 0.12E-6
+LD    = 0.35E-6
+DELTA = 0.25
+THETA = 0.060
+ETA   = 0.030
+KAPPA = 0.0
+WD    = -0.5E-6

***********************************************
*          SLOW P-Channel transistor          *
*           UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family        *
*                10-Jan.-1995                 *
***********************************************
.Model MHCPES PMOS
+LEVEL = 3
+KP    = 19.6E-6
+VTO   = -0.91
+TOX   = 54.0E-9
+NSUB  = 3.0E16
+GAMMA = 1.02
+PHI   = 0.65
+VMAX  = 190E4
+RS    = 100
+RD    = 100
+XJ    = 0.65E-6
+LD    = 0.10E-6
+DELTA = 2.35
+THETA = 0.120
+ETA   = 0.380
+KAPPA = 0.0
+WD    = -0.5E-6


.MODEL  INT D

****************************************
*   START OF SUB-CIRCUIT DESCRIPTION   *
*            MARCH 28, 1995            *
****************************************


*****SLOW.CIR*****

****Version 1.04 Added Inverter****
.SUBCKT INV4S   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPES W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2 60 60  MHCNES W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
.ENDS


.SUBCKT INP0S  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  3  100
MP1 3 50 50 50  MHCPES W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 3 60 60 60  MHCNES W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
.ENDS

.SUBCKT INP1S  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNES W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
MP2 3  4 50 50  MHCPES W=88U L=2.4U AD=290P AS=550P PD=10U PS=100U
MN2 3  4 60 60  MHCNES W=56U L=2.4U AD=162P AS=550P PD=10U PS= 75U
.ENDS

.SUBCKT INP1TS  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W= 20U L=2.4U AD=100P AS=100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNES W= 35U L=2.4U AD=260P AS=260P PD= 70U PS= 20U
MP2 3  4  5 50  MHCPES W= 88U L=2.4U AD=290P AS=550P PD=107U PS=195U
MN2 3  4 60 60  MHCNES W= 56U L=2.4U AD=162P AS=550P PD= 55U PS=162U
D1 50  5  INT
MP4 3  6 50 50  MHCPES W=6.4U L=4.0U AD= 60P AS= 60P PD= 13U PS= 24U
MN4 3  4 60 60  MHCNES W=185U L=2.4U AD=740P AS=740P PD= 50U PS=185U
MP5 6  3 50 50  MHCPES W=6.4U L=3.2U AD= 50P AS= 50P PD= 10U PS= 20U
MN5 6  3 60 60  MHCNES W=6.4U L=3.2U AD= 50P AS= 50P PD= 10U PS= 20U
.ENDS

.SUBCKT INP2S  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W= 20U L=2.4U AD= 100P AS=100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNES W= 35U L=2.4U AD= 260P AS=260P PD= 70U PS= 20U
MP2 3  4 50 50  MHCPES W=176U L=2.4U AD= 580P AS=580P PD=10U PS=200U
MN2 3  4 60 60  MHCNES W=112U L=2.4U AD= 325P AS=580P PD=10U PS=150U
.ENDS

.SUBCKT INP2TS  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W= 20U L=2.4U AD= 100P AS= 100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNES W= 35U L=2.4U AD= 260P AS= 260P PD= 70U PS= 20U
MP2 3  4  5 50  MHCPES W=176U L=2.4U AD= 580P AS=1100P PD=215U PS=390U
MN2 3  4 60 60  MHCNES W=440U L=2.4U AD=1320P AS=1840P PD=190U PS=650U
D1 50  5   INT
MP4 3  6 50 50  MHCPES W=6.4U L=4.0U AD=  60P AS=  60P PD= 13U PS= 24U
MP5 6  3 50 50  MHCPES W=6.4U L=3.2U AD=  50P AS=  50P PD= 10U PS= 20U
MN5 6  3 60 60  MHCNES W=6.4U L=3.2U AD=  50P AS=  50P PD= 10U PS= 20U
.ENDS


.SUBCKT SMT1S  2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HC14 CMOS INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W=20U L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNES W=35U L=2.4U AD=140P AS=140P PD=50U PS=35U
MP2 5  4 50 50  MHCPES W=36U L=2.4U AD=140P AS=140P PD=50U PS=35U
MN2 6  4 60 60  MHCNES W=16U L=2.4U AD= 70P AS= 70P PD=15U PS=17U
MP3 3  4  5 50  MHCPES W=44U L=2.4U AD=220P AS=220P PD=60U PS=44U
MN3 3  4  6  6  MHCNES W=17U L=2.4U AD= 70P AS= 70P PD=15U PS=16U
MP4 5  3 60 50  MHCPES W=36U L=2.4U AD=150P AS=150P PD=60U PS=36U
MN4 6  3 50  6  MHCNES W= 6U L=  4U AD= 25P AS= 25P PD=10U PS= 6U
.ENDS


.SUBCKT SMTTL1S  2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HCT14 WITH TTL INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPES W= 20U L=2.4U AD= 100P AS= 100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNES W= 35U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
D1  50  7  INT
MP2 5  4  7  7  MHCPES W= 36U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
MN2 6  4 60 60  MHCNES W=216U L=2.4U AD= 860P AS= 860P PD=140U PS=216U
MP3 3  4  5 50  MHCPES W= 54U L=2.4U AD= 220P AS= 220P PD= 60U PS= 44U
MN3 3  4  6  6  MHCNES W=257U L=2.4U AD=1000P AS=1000P PD=150U PS=257U
MP4 5  3 60 50  MHCPES W= 32U L=  4U AD= 120P AS= 120P PD=100U PS= 32U
MN4 6  3 50  6  MHCNES W= 14U L=  4U AD= 100P AS= 100P PD= 30U PS= 24U
MP5 8  3 50 50  MHCPES W= 10U L=2.4U AD=  40P AS=  40P PD= 16U PS= 10U
MN5 8  3 60 60  MHCNES W=  5U L=2.4U AD=  20P AS=  20P PD= 12U PS=  5U
MP6 3  8 50 50  MHCPES W=  6U L=8.0U AD=  30P AS=  30P PD= 16U PS=  6U
.ENDS


.SUBCKT INVS   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPES W=364U L=2.4U AD=500P  AS=500P PD=10U PS=430U
MN1 3  2 60 60  MHCNES W=184U L=2.4U AD=275P  AS=275P PD=10U PS=270U
.ENDS


.SUBCKT NANDS  2  3  4  50  60
*INTERNAL NAND
*IN1 = 2, IN2 = 3, OUT = 4, VCC= 50, GND = 60
MP1 4  2  50  50  MHCPES W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MP2 4  3  50  50  MHCPES W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MN1 4  2   5  60  MHCNES W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
MN2 5  3  60  60  MHCNES W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
.ENDS


.SUBCKT LLCS  2  3  40  50  60
* LEVEL CONVERTER
* INA = 2,  OUT = 3,  VEE = 40,  VCC = 50,  GND =  60
MP4 4  2  50  50  MHCPES W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN4 4  2  60  60  MHCNES W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
MP1 5  4  50  50  MHCPES W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MP2 6  2  50  50  MHCPES W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MN1 5  6  40  40  MHCNES W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MN2 6  5  40  40  MHCNES W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MP3 7  6  50  50  MHCPES W= 10U  L= 4.0U AD= 40P AS= 40P PD= 20U PS= 10U
MN3 7  6  40  40  MHCNES W=  5U  L= 4.0U AD= 20P AS= 20P PD= 10U PS=  5U
MP5 3  7  50  50  MHCPES W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN5 3  7  40  40  MHCNES W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
.ENDS

.SUBCKT SWITCH1S  2  8  9  40  50
* ANALOG SWITCH
* INPUT = 2   Y = 8  Z = 9  VEE = 40  VCC =50
MP1 3  2  50  50  MHCPES W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNES W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPES W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNES W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 8  4   5  50  MHCPES W= 216U L=2.4U AD= 900P AS= 900P PD=100U PS= 216U
MN5 8  3   5   5  MHCNES W= 108U L=2.4U AD= 430P AS= 430P PD= 50U PS= 108U
MN6 5  4  40  40  MHCNES W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  4   8  50  MHCPES W=1068U L=2.4U AD=2500P AS=2500P PD= 10U PS=1068U
MN7 9  3   8   5  MHCNES W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS

.SUBCKT SWITCH2S  2  8  9  50  60
* ANALOG SWITCH
* INPUT= 2   Y= 8   Z= 9  VCC= 50   GND= 60
MP1 3  2  50  50  MHCPES W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  60  60  MHCNES W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPES W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  60  60  MHCNES W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 5  3   8  50  MHCPES W=  85U L=2.4U AD= 355P AS= 355P PD= 40U PS=  85U
MN5 5  4   8   5  MHCNES W=  42U L=2.4U AD= 170P AS= 170P PD= 20U PS=  42U
MN6 5  3  60  60  MHCNES W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  3   8  50  MHCPES W=1900U L=2.4U AD=2500P AS=2500P PD= 10U PS=1900U
MN7 9  4   8   5  MHCNES W= 576U L=2.4U AD=1200P AS=1200P PD= 10U PS= 576U
.ENDS

.SUBCKT SWITCH3S  2  8  9  40  50
* ANALOG SWITCH
* INPUT = 2   Y = 8  Z = 9  VEE = 40  VCC = 50
MP1 3  2  50  50  MHCPES W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNES W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPES W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNES W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 9  3   8  50  MHCPES W=1168U L=2.4U AD=2730P AS=2730P PD= 10U PS=1168U
MN5 9  4   8  40  MHCNES W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS


.SUBCKT BUSOUTPS  2   3   4   50   60
* INPUT = 2  OEN = 3 (LOW)  OUT = 4  VCC = 50  GND = 60
* 3-STATE BUS OUTPUT
MP1 5  3   50  50  MHCPES W= 90U  L=2.4U AD= 360P AS= 360P PD= 30U PS=360U
MN1 5  3   60  60  MHCNES W= 40U  L=2.4U AD= 160P AS= 160P PD= 20U PS= 40U
MP2 6  2   50  50  MHCPES W=480U  L=2.4U AD=1800P AS=1800P PD=100U PS=480U
MN2 7  2   60  60  MHCNES W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MP3 7  3    6  50  MHCPES W=280U  L=2.4U AD=1120P AS=1120P PD= 55U PS=280U
MN3 7  3   60  60  MHCNES W=160U  L=2.4U AD= 640P AS= 640P PD= 40U PS=160U
MP4 6  5   50  50  MHCPES W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MN4 7  5    7  60  MHCNES W=190U  L=2.4U AD= 760P AS= 760P PD= 45U PS=190U
R1  6  8  200
R2  7  9  200
MP5 4  8   50  50  MHCPES W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN5 4  9   60  60  MHCNES W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R3  8  10 100
R4  9  11 100
MP6 4  10  50  50  MHCPES W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN6 4  11  60  60  MHCNES W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R5 10  12  50
R6 11  13  50
MP7 4  12  50  50  MHCPES W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN7 4  13  60  60  MHCNES W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
.ENDS


.SUBCKT OUTUS  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPES W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN1 3 4 60 60  MHCNES W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPES W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN2 3 5 60 60  MHCNES W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPES W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN3 3 6 60 60  MHCNES W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
.ENDS

.SUBCKT OUTPS  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPES W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN1 3 4 60 60  MHCNES W=140U L=2.4U AD=200P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPES W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN2 3 5 60 60  MHCNES W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPES W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN3 3 6 60 60  MHCNES W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
.ENDS

*******************************************************************
*******************************************************************

******CIR_SLOW_HC TYPES******


.SUBCKT INV0  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP0S
XOUTP 25  30  50  60    OUTUS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  30   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV1  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1S
XINV  25  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV2  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP2S
XINV  25  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INVSMT  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    SMT1S
XINV  25  30  50  60    INVS
XOUTP 30  40  50  60    OUTPS
L1  80  50   3.54NH
L2  60  90   3.54NH
L3   2  20   3.54NH
L4  40   3   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NINV1  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1S
XINV0 25  30  50  60    INVS
XINV1 30  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NANDINV 2  5  3  80  90
*INVERTING 2-NAND
*EN = 5, IN = 2, OUT = 3, VCC = 80, GND = 90
XIN1  20  25      50  60   INP2S
XIN2  30  35      50  60   INP2S
XNAND 25  35  36  50  60   NANDS
XOUT  36  40      50  60   OUTPS
L1     2  20   4.28NH
L2     5  30   4.28NH
L3    40   3   6.08NH
L4    80  50   6.08NH
L5    60  90   6.08NH
C1    20  90   1.5P
C2    30  90   1.5P
C3    40  90   1.5P
C4    50  90   1.5P
C5    60  90   1.5P
.ENDS


.SUBCKT SWI1  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP2S
XLC  25  30  40  50  60  LLCS
XAS  30   3   4  40  50  SWITCH1S
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS



.SUBCKT SWI2  2  3  4  80  90
* INP = 2  Y = 3  Z = 4  VCC = 80  GND = 90
*XINP  20  25  50  60      INP2S
****Version 1.04 Inserted inverter****
XINP  20  250  50  60      INP2S
XINV  250  25  50  60      INV4S
XAS   25   8   9  50  60  SWITCH2S
L1  80  50   3.53NH
L2  60  90   3.54NH
L3   2  20   3.53NH
L4   8   3   3.54NH
L5   9   4   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
C5  4   90   1.5P
.ENDS


.SUBCKT SWI3  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP1S
XLC  25  30  40  50  60  LLCS
XAS  30   3   4  40  50  SWITCH3S
L1  80  50   5.97NH
L2  70  40   5.97NH
L3  60  90   5.97NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT NINV3  2  5  3  80  90
* INP = 2  OEN = 5(LOW)  OUT = 3   VCC = 80  GND = 90
XINP      20  25  50  60      INP2S
XINV      25  30  50  60      INVS
XBUSOUTP  30  15  35  50  60  BUSOUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   6.87NH
L4   5  15   5.97NH
L5  35   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C4  20  90   1.5P
C5  15  90   1.5P
C6   3  90   1.5P
.ENDS



******CIR_SLOW_HCT TYPES******

.SUBCKT INV0T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP0S
XOUTP 25  30  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  30   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV1T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1TS
XINV  25  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV2T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP2TS
XINV  25  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INVSMTT  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    SMTTL1S
XINV  25  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   3.54NH
L2  60  90   3.54NH
L3   2  20   3.54NH
L4  40   3   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NINV1T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1TS
XINV0 25  30  50  60    INVS
XINV1 30  35  50  60    INVS
XOUTP 35  40  50  60    OUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NANDINVT 2  5  3  80  90
*INVERTING 2-NAND
*EN = 5, IN = 2, OUT = 3, VCC = 80, GND = 90
XIN1  20  25      50  60   INP2TS
XIN2  30  35      50  60   INP2TS
XNAND 25  35  36  50  60   NANDS
XOUT  36  40      50  60   OUTPS
L1     2  20   5.29NH
L2     5  30   4.28NH
L3    40   3   3.78NH
L4    80  50   6.08NH
L5    60  90   6.08NH
C1    20  90   1.5P
C2    30  90   1.5P
C3    40  90   1.5P
C4    50  90   1.5P
C5    60  90   1.5P
.ENDS


.SUBCKT SWI1T  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP2TS
XLC  25  30  40  50  60  LLCS
XAS  30   3   4  40  50  SWITCH1S
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT SWI2T  2  3  4  80  90
* INP = 2  Y = 3  Z = 4  VCC = 80  GND = 90
*XINP  20  25  50  60      INP1TS
****Version 1.04 Inserted inverter****
XINP  20  250  50  60      INP1TS
XINV  250  25  50  60      INV4S
XAS   25   8   9  50  60  SWITCH2S
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4   8   3   5.97NH
L5   9   4   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
C5  4   90   1.5P
.ENDS


.SUBCKT SWI3T  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP1TS
XLC  25  30  40  50  60  LLCS
XAS  30   3   4  40  50  SWITCH3S
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT NINV3T  2  5  3  80  90
*
* INP = 2  OEN = 5(LOW)  OUT = 3   VCC = 80  GND = 90
XINP      20  25  50  60      INP2TS
XINV      25  30  50  60      INVS
XBUSOUTP  30  15  35  50  60  BUSOUTPS
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   6.87NH
L4   5  15   5.97NH
L5  35   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C4  20  90   1.5P
C5  15  90   1.5P
C6   3  90   1.5P
.ENDS


***********************************************************
