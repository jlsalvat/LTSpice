* HCMOS Subcircuit and Primitive Elements Library
* HC_TNOMI.CIR
* Nominal Process Corner
* Standard Logic Product Group
* Philips Semiconductors
*
* Version Date       By   Remarks
* ---------------------------------------------------------------------
*    1.05 10/27/2005 RRV  Updated HC/T04 and HCU04 models
*    1.04 09/22/2003 RM   Active High Enable for SWI2 and SWI2T
*
************************************************
*         NOMINAL N-Channel Transistor         *
*            UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family         *
*                10-Jan.-1995                  *
************************************************
.Model MHCNEN NMOS
+LEVEL = 3
+KP    = 45.3E-6
+VTO   = 0.72
+TOX   = 51.5E-9
+NSUB  = 2.8E15
+GAMMA = 0.94
+PHI   = 0.65
+VMAX  = 150E3
+RS    = 40
+RD    = 40
+XJ    = 0.11E-6
+LD    = 0.52E-6
+DELTA = 0.315
+THETA = 0.054
+ETA   = 0.025
+KAPPA = 0.0
+WD    = 0.0

***********************************************
*        NOMINAL P-Channel transistor         *
*           UCB-3 Parameter Set               *
*         HIGH-SPEED CMOS Logic Family        *
*               10-Jan.-1995                  *
***********************************************
.Model MHCPEN PMOS
+LEVEL = 3
+KP    = 22.1E-6
+VTO   = -0.71
+TOX   = 51.5E-9
+NSUB  = 3.3E16
+GAMMA = 0.92
+PHI   = 0.65
+VMAX  = 970E3
+RS    = 80
+RD    = 80
+XJ    = 0.63E-6
+LD    = 0.23E-6
+DELTA = 2.24
+THETA = 0.108
+ETA   = 0.322
+KAPPA = 0.0
+WD    = 0.0


.MODEL  INT D


****************************************
*   START OF SUB-CIRCUIT DESCRIPTION   *
*            MARCH 28, 1995            *
****************************************

*****NOMIN.CIR*****

****Version 1.04 Added Inverter****
.SUBCKT INV4N   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPEN W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2 60 60  MHCNEN W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
.ENDS


.SUBCKT INP0N  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  3  100
MP1 3 50 50 50  MHCPEN W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 3 60 60 60  MHCNEN W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
.ENDS

.SUBCKT INP1N  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W=20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEN W=35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
MP2 3  4 50 50  MHCPEN W=88U L=2.4U AD=290P AS=550P PD=10U PS=100U
MN2 3  4 60 60  MHCNEN W=56U L=2.4U AD=162P AS=550P PD=10U PS= 75U
.ENDS

.SUBCKT INP1TN  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W= 20U L=2.4U AD=100P AS=100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNEN W= 35U L=2.4U AD=260P AS=260P PD= 70U PS= 20U
MP2 3  4  5 50  MHCPEN W= 88U L=2.4U AD=290P AS=550P PD=107U PS=195U
MN2 3  4 60 60  MHCNEN W= 56U L=2.4U AD=162P AS=550P PD= 55U PS=162U
D1 50  5  INT
MP4 3  6 50 50  MHCPEN W=6.4U L=4.0U AD= 60P AS= 60P PD=13U PS= 24U
MN4 3  4 60 60  MHCNEN W=185U L=2.4U AD=740P AS=740P PD=50U PS=185U
MP5 6  3 50 50  MHCPEN W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
MN5 6  3 60 60  MHCNEN W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
.ENDS

.SUBCKT INP2N  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W= 20U L=2.4U AD=100P AS=100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEN W= 35U L=2.4U AD=260P AS=260P PD=70U PS= 20U
MP2 3  4 50 50  MHCPEN W=176U L=2.4U AD=580P AS=580P PD=10U PS=200U
MN2 3  4 60 60  MHCNEN W=112U L=2.4U AD=325P AS=580P PD=10U PS=150U
.ENDS

.SUBCKT INP2TN  2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W= 20U L=2.4U AD=100P AS= 100P PD=40U PS= 20U
MN1 4 60 60 60  MHCNEN W= 35U L=2.4U AD=260P AS= 260P PD=70U PS= 20U
MP2 3  4  5 50  MHCPEN W=176U L=2.4U AD=580P AS=1100P PD=10U PS=200U
MN2 3  4 60 60  MHCNEN W=112U L=2.4U AD=325P AS=1100P PD=10U PS=150U
D1 50  5   INT
MP4 3  6 50 50  MHCPEN W=6.4U L=4.0U AD= 60P AS= 60P PD=13U PS= 24U
MN4 3  4 60 60  MHCNEN W=348U L=2.4U AD=740P AS=740P PD=50U PS=348U
MP5 6  3 50 50  MHCPEN W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
MN5 6  3 60 60  MHCNEN W=6.4U L=3.2U AD= 50P AS= 50P PD=10U PS= 20U
.ENDS


.SUBCKT SMT1N  2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HC14 CMOS INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W=20U L=2.4U AD=100P AS=100P PD=40U PS=20U
MN1 4 60 60 60  MHCNEN W=35U L=2.4U AD=140P AS=140P PD=50U PS=35U
MP2 5  4 50 50  MHCPEN W=36U L=2.4U AD=140P AS=140P PD=50U PS=35U
MN2 6  4 60 60  MHCNEN W=16U L=2.4U AD= 70P AS= 70P PD=15U PS=17U
MP3 3  4  5 50  MHCPEN W=44U L=2.4U AD=220P AS=220P PD=60U PS=44U
MN3 3  4  6  6  MHCNEN W=17U L=2.4U AD= 70P AS= 70P PD=15U PS=16U
MP4 5  3 60 50  MHCPEN W=36U L=2.4U AD=150P AS=150P PD=60U PS=36U
MN4 6  3 50  6  MHCNEN W= 6U L=  4U AD= 25P AS= 25P PD=10U PS= 6U
.ENDS


.SUBCKT SMTTL1N  2  3  50  60
* SCHMITT-TRIGGER INPUT FOR HCT14 WITH TTL INPUT LEVELS
*IN=2, OUT=3, VCC=50, GND=60
R1  2  4  100
MP1 4 50 50 50  MHCPEN W= 20U L=2.4U AD= 100P AS= 100P PD= 40U PS= 20U
MN1 4 60 60 60  MHCNEN W= 35U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
D1  50  7  INT
MP2 5  4  7  7  MHCPEN W= 36U L=2.4U AD= 140P AS= 140P PD= 50U PS= 35U
MN2 6  4 60 60  MHCNEN W=216U L=2.4U AD= 860P AS= 860P PD=140U PS=216U
MP3 3  4  5 50  MHCPEN W= 54U L=2.4U AD= 220P AS= 220P PD= 60U PS= 44U
MN3 3  4  6  6  MHCNEN W=257U L=2.4U AD=1000P AS=1000P PD=150U PS=257U
MP4 5  3 60 50  MHCPEN W= 32U L=  4U AD= 120P AS= 120P PD=100U PS= 32U
MN4 6  3 50  6  MHCNEN W= 14U L=  4U AD= 100P AS= 100P PD= 30U PS= 24U
MP5 8  3 50 50  MHCPEN W= 10U L=2.4U AD=  40P AS=  40P PD= 16U PS= 10U
MN5 8  3 60 60  MHCNEN W=  5U L=2.4U AD=  20P AS=  20P PD= 12U PS=  5U
MP6 3  8 50 50  MHCPEN W=  6U L=8.0U AD=  30P AS=  30P PD= 16U PS=  6U
.ENDS


.SUBCKT INVN   2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
MP1 3  2 50 50  MHCPEN W=364U L=2.4U AD=500P  AS=500P PD=10U PS=430U
MN1 3  2 60 60  MHCNEN W=184U L=2.4U AD=275P  AS=275P PD=10U PS=270U
.ENDS


.SUBCKT NANDN  2  3  4  50  60
*INTERNAL NAND
*IN1 = 2, IN2 = 3, OUT = 4, VCC= 50, GND = 60
MP1 4  2  50  50  MHCPEN W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MP2 4  3  50  50  MHCPEN W=112U  L=2.4U AD=150P AS=300P PD= 75U PS=150U
MN1 4  2   5  60  MHCNEN W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
MN2 5  3  60  60  MHCNEN W=300U  L=2.4U AD=300P AS=300P PD=300U PS=300U
.ENDS


.SUBCKT LLCN  2  3  40  50  60
* LEVEL CONVERTER
* INA = 2,  OUT = 3,  VEE = 40,  VCC = 50,  GND =  60
MP4 4  2  50  50  MHCPEN W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN4 4  2  60  60  MHCNEN W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
MP1 5  4  50  50  MHCPEN W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MP2 6  2  50  50  MHCPEN W=135U  L= 2.4U AD=500P AS=500P PD=100U PS=135U
MN1 5  6  40  40  MHCNEN W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MN2 6  5  40  40  MHCNEN W=6.4U  L=18.8U AD= 25P AS= 25P PD= 20U PS=6.4U
MP3 7  6  50  50  MHCPEN W= 10U  L= 4.0U AD= 40P AS= 40P PD= 20U PS= 10U
MN3 7  6  40  40  MHCNEN W=  5U  L= 4.0U AD= 20P AS= 20P PD= 10U PS=  5U
MP5 3  7  50  50  MHCPEN W= 30U  L= 2.4U AD=120P AS=120P PD= 40U PS= 30U
MN5 3  7  40  40  MHCNEN W= 15U  L= 2.4U AD= 60P AS= 60P PD= 20U PS= 15U
.ENDS

.SUBCKT SWITCH1N  2  8  9  40  50
* ANALOG SWITCH
* INPUT = 2,   Y = 8,  Z = 9,  VEE = 40,  VCC =50
MP1 3  2  50  50  MHCPEN W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNEN W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEN W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNEN W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 8  4   5  50  MHCPEN W= 216U L=2.4U AD= 900P AS= 900P PD=100U PS= 216U
MN5 8  3   5   5  MHCNEN W= 108U L=2.4U AD= 430P AS= 430P PD= 50U PS= 108U
MN6 5  4  40  40  MHCNEN W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  4   8  50  MHCPEN W=1068U L=2.4U AD=2500P AS=2500P PD= 10U PS=1068U
MN7 9  3   8   5  MHCNEN W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS

.SUBCKT SWITCH2N  2  8  9  50  60
* ANALOG SWITCH
* INPUT= 2   Y= 8   Z= 9  VCC= 50   GND= 60
MP1 3  2  50  50  MHCPEN W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  60  60  MHCNEN W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEN W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  60  60  MHCNEN W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 5  3   8  50  MHCPEN W=  85U L=2.4U AD= 355P AS= 355P PD= 40U PS=  85U
MN5 5  4   8   5  MHCNEN W=  42U L=2.4U AD= 170P AS= 170P PD= 20U PS=  42U
MN6 5  3  60  60  MHCNEN W= 145U L=2.4U AD= 600P AS= 600P PD= 75U PS= 145U
MP7 9  3   8  50  MHCPEN W=1900U L=2.4U AD=2500P AS=2500P PD= 10U PS=1900U
MN7 9  4   8   5  MHCNEN W= 576U L=2.4U AD=1200P AS=1200P PD= 10U PS= 576U
.ENDS

.SUBCKT SWITCH3  2  8  9  40  50
* ANALOG SWITCHN
* INPUT = 2   Y = 8  Z = 9  VEE = 40  VCC = 50
MP1 3  2  50  50  MHCPEN W=  88U L=2.4U AD= 350P AS= 350P PD=100U PS=  88U
MN1 3  2  40  40  MHCNEN W=  56U L=2.4U AD= 225P AS= 225P PD= 70U PS=  56U
MP4 4  3  50  50  MHCPEN W= 350U L=2.4U AD= 900P AS= 900P PD=200U PS= 350U
MN4 4  3  40  40  MHCNEN W= 150U L=2.4U AD= 400P AS= 400P PD=100U PS= 150U
MP5 9  3   8  50  MHCPEN W=1168U L=2.4U AD=2730P AS=2730P PD= 10U PS=1168U
MN5 9  4   8  40  MHCNEN W= 312U L=2.4U AD=1200P AS=1200P PD= 10U PS= 312U
.ENDS


.SUBCKT BUSOUTPN  2   3   4   50   60
* INPUT = 2  OEN = 3 (LOW)  OUT = 4  VCC = 50  GND = 60
* 3-STATE BUS OUTPUT
MP1 5  3   50  50  MHCPEN W= 90U  L=2.4U AD= 360P AS= 360P PD= 30U PS=360U
MN1 5  3   60  60  MHCNEN W= 40U  L=2.4U AD= 160P AS= 160P PD= 20U PS= 40U
MP2 6  2   50  50  MHCPEN W=480U  L=2.4U AD=1800P AS=1800P PD=100U PS=480U
MN2 7  2   60  60  MHCNEN W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MP3 7  3    6  50  MHCPEN W=280U  L=2.4U AD=1120P AS=1120P PD= 55U PS=280U
MN3 7  3   60  60  MHCNEN W=160U  L=2.4U AD= 640P AS= 640P PD= 40U PS=160U
MP4 6  5   50  50  MHCPEN W=240U  L=2.4U AD=1000P AS=1000P PD= 50U PS=240U
MN4 7  5    7  60  MHCNEN W=190U  L=2.4U AD= 760P AS= 760P PD= 45U PS=190U
R1  6  8  200
R2  7  9  200
MP5 4  8   50  50  MHCPEN W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN5 4  9   60  60  MHCNEN W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R3  8  10 100
R4  9  11 100
MP6 4  10  50  50  MHCPEN W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN6 4  11  60  60  MHCNEN W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
R5 10  12  50
R6 11  13  50
MP7 4  12  50  50  MHCPEN W=540U  L=2.4U AD=1500P AS=1500P PD=10U PS=540U
MN7 4  13  60  60  MHCNEN W=233U  L=2.4U AD= 750P AS= 750P PD=10U PS=233U
.ENDS

.SUBCKT OUTUN 2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPEN W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN1 3 4 60 60  MHCNEN W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPEN W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN2 3 5 60 60  MHCNEN W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPEN W=485U L=2.4U AD=1200P AS=530P PD=10U PS=180U
MN3 3 6 60 60  MHCNEN W=222U L=2.4U AD=530P AS=300P PD=10U PS=130U
.ENDS

.SUBCKT OUTPN 2  3  50  60
*IN=2, OUT=3, VCC=50, GND=60
R1  2 4 100
MP1 3 4 50 50  MHCPEN W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN1 3 4 60 60  MHCNEN W=140U L=2.4U AD=200P AS=300P PD=10U PS=130U
R2  4 5 50
MP2 3 5 50 50  MHCPEN W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN2 3 5 60 60  MHCNEN W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
R3  5 6 50
MP3 3 6 50 50  MHCPEN W=360U L=2.4U AD=400P AS=400P PD=10U PS=180U
MN3 3 6 60 60  MHCNEN W=140U L=2.4U AD=200P AS=200P PD=10U PS=130U
.ENDS

*******************************************************************
*******************************************************************

******CIR_NOMIN-HC TYPES******

.SUBCKT INV0  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP0N
XOUTP 25  30  50  60    OUTUN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  30   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV1  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1N
XINV  25  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV2  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP2N
XINV  25  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INVSMT  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    SMT1N
XINV  25  30  50  60    INVN
XOUTP 30  40  50  60    OUTPN
L1  80  50   3.54NH
L2  60  90   3.54NH
L3   2  20   3.54NH
L4  40   3   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NINV1  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1N
XINV0 25  30  50  60    INVN
XINV1 30  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NANDINV 2  5  3  80  90
*INVERTING 2-NAND
*EN = 5, IN = 2, OUT = 3, VCC = 80, GND = 90
XIN1  20  25      50  60   INP2N
XIN2  30  35      50  60   INP2N
XNAND 25  35  36  50  60   NANDN
XOUT  36  40      50  60   OUTPN
L1     2  20   4.28NH
L2     5  30   4.28NH
L3    40   3   6.08NH
L4    80  50   6.08NH
L5    60  90   6.08NH
C1    20  90   1.5P
C2    30  90   1.5P
C3    40  90   1.5P
C4    50  90   1.5P
C5    60  90   1.5P
.ENDS


.SUBCKT SWI1  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP2N
XLC  25  30  40  50  60  LLCN
XAS  30   3   4  40  50  SWITCH1N
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT SWI2  2  3  4  80  90
* INP = 2  Y = 3  Z = 4  VCC = 80  GND = 90
*XINP  20  25  50  60      INP2N
****Version 1.04 Inserted inverter****
XINP  20  250  50  60      INP2N
XINV  250  25  50  60      INV4N
XAS   25   8   9  50  60  SWITCH2N
L1  80  50   3.53NH
L2  60  90   3.54NH
L3   2  20   3.53NH
L4   8   3   3.54NH
L5   9   4   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
C5  4   90   1.5P
.ENDS


.SUBCKT SWI3  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP1N
XLC  25  30  40  50  60  LLCN
XAS  30   3   4  40  50  SWITCH3N
L1  80  50   5.97NH
L2  70  40   5.97NH
L3  60  90   5.97NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT NINV3  2  5  3  80  90
* INP = 2  OEN = 5(LOW)  OUT = 3   VCC = 80  GND = 90
XINP      20  25  50  60      INP2N
XINV      25  30  50  60      INVN
XBUSOUTP  30  15  35  50  60  BUSOUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   6.87NH
L4   5  15   5.97NH
L5  35   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C4  20  90   1.5P
C5  15  90   1.5P
C6   3  90   1.5P
.ENDS



******CIR_NOMIN-HCT TYPES******

.SUBCKT INV0T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP0N
XOUTP 25  30  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  30   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV1T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1TN
XINV  25  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INV2T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP2TN
XINV  25  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT INVSMTT  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    SMTTL1N
XINV  25  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   3.54NH
L2  60  90   3.54NH
L3   2  20   3.54NH
L4  40   3   3.54NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NINV1T  2  3  80 90
*IN=2, OUT=3, VCC=80, GND=90
XINP  20  25  50  60    INP1TN
XINV0 25  30  50  60    INVN
XINV1 30  35  50  60    INVN
XOUTP 35  40  50  60    OUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4  40   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
.ENDS


.SUBCKT NANDINVT 2  5  3  80  90
*INVERTING 2-NAND
*EN = 5, IN = 2, OUT = 3, VCC = 80, GND = 90
XIN1  20  25      50  60   INP2TN
XIN2  30  35      50  60   INP2TN
XNAND 25  35  36  50  60   NANDN
XOUT  36  40      50  60   OUTPN
L1     2  20   5.29NH
L2     5  30   4.28NH
L3    40   3   3.78NH
L4    80  50   6.08NH
L5    60  90   6.08NH
C1    20  90   1.5P
C2    30  90   1.5P
C3    40  90   1.5P
C4    50  90   1.5P
C5    60  90   1.5P
.ENDS


.SUBCKT SWI1T  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP2TN
XLC  25  30  40  50  60  LLCN
XAS  30   3   4  40  50  SWITCH1N
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT SWI2T  2  3  4  80  90
* INP = 2  Y = 3  Z = 4  VCC = 80  GND = 90
*XINP  20  25  50  60      INP1TN
****Version 1.04 Inserted inverter****
XINP  20  250  50  60      INP1TN
XINV  250  25  50  60      INV4N
XAS   25   8   9  50  60  SWITCH2N
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   5.97NH
L4   8   3   5.97NH
L5   9   4   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C3  20  90   1.5P
C4  3   90   1.5P
C5  4   90   1.5P
.ENDS


.SUBCKT SWI3T  2  3  4  70  80  90
* INP = 2  Y = 3  Z = 4  VEE = 70  VCC = 80  GND = 90
XINP 20  25  50  60      INP1TN
XLC  25  30  40  50  60  LLCN
XAS  30   3   4  40  50  SWITCH3N
L1  80  50   6.08NH
L2  70  40   6.08NH
L3  60  90   6.08NH
L4   2  20   4.28NH
C1  50  90   1.5P
C2  40  90   1.5P
C3  60  90   1.5P
C4  20  90   1.5P
C5  3   90   1.5P
C6  4   90   1.5P
.ENDS


.SUBCKT NINV3T  2  5  3  80  90
*
* INP = 2  OEN = 5(LOW)  OUT = 3   VCC = 80  GND = 90
XINP      20  25  50  60      INP2TN
XINV      25  30  50  60      INVN
XBUSOUTP  30  15  35  50  60  BUSOUTPN
L1  80  50   6.87NH
L2  60  90   6.87NH
L3   2  20   6.87NH
L4   5  15   5.97NH
L5  35   3   5.97NH
C1  50  90   1.5P
C2  60  90   1.5P
C4  20  90   1.5P
C5  15  90   1.5P
C6   3  90   1.5P
.ENDS


***********************************************************
